module AHBDVP(

);



endmodule